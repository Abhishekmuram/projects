class mon extends uvm_monitor;
`uvm_component_utils(mon)

transaction tr;
virtual sram_if sif;
uvm_analysis_port#(transaction)send;

function new(string name="mon",uvm_component parent=null);
super.new(name,parent);
endfunction


virtual function void build_phase(uvm_phase phase);
super.build_phase(phase);
tr=transaction::type_id::create("tr");
send=new("send",this);
if(!uvm_config_db #(virtual sram_if)::get(this,"","sif",sif))
`uvm_error(get_type_name(),"unable to access interface");
endfunction

virtual task run_phase(uvm_phase phase);
    forever begin
      repeat(2) @(posedge sif.clk);
    tr.wr_enable=sif.wr_enable;
    tr.addr=sif.addr;
    tr.din=sif.din;
    tr.dout=sif.dout;
     `uvm_info("mon",$sformatf("wr_enable:%0b addr:%0d din:%0d dout:%0d",tr.wr_enable,tr.addr,tr.din,tr.dout),UVM_NONE);
        send.write(tr);
    end
   endtask 
 
endclass

