interface mux_if();

logic a;
logic b;
logic s;
logic y;

endinterface

