class test extends uvm_test;
`uvm_component_utils(test)

function new(string name="test",uvm_component parent=null);
super.new(name,parent);
endfunction

env e;
//write_data wd;
//read_data  rd;
write_read  wr;
//write_err  er;



virtual function void build_phase(uvm_phase phase);
super.build_phase(phase);
e=env::type_id::create("e",this);
//wd=write_data::type_id::create("wd");
//rd=read_data::type_id::create("rd");
wr=write_read::type_id::create("wr");
//er=write_err::type_id::create("er");
endfunction

virtual task run_phase(uvm_phase phase);
phase.raise_objection(this);

wr.start(e.a.seqr);

#20;

phase.drop_objection(this);
endtask
endclass




