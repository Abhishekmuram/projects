interface and_if();
  logic a;
  logic b;
  logic y;
endinterface
