interface sram_if();

logic clk,rst;
logic wr_enable;
logic [4:0]addr;
logic [4:0]din;
logic [4:0]dout;


endinterface
