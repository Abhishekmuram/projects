import uvm_pkg::*;
`include "uvm_macros.svh"
`include "dut.sv"
`include "interface.sv"
`include "sequence_item.sv"
`include "sequencer.sv"
//`include "seq_1.sv"
//`include "seq_2.sv"
`include "seq_3.sv"
//`include "seq_4.sv"
`include "driver.sv"
`include "monitor.sv"
`include "agent.sv"
`include "sco.sv"

`include "env.sv"
`include "test.sv"
//`include "top.sv"


module tb;
  
  
  apb_if aif();
  
  apb_ram dut (.presetn(aif.presetn), .pclk(aif.pclk), .psel(aif.psel), .penable(aif.penable), .pwrite(aif.pwrite), .paddr(aif.paddr), .pwdata(aif.pwdata), .prdata(aif.prdata), .pready(aif.pready), .pslverr(aif.pslverr));
  
  initial begin
    aif.pclk = 0;
  end
 
   always #10 aif.pclk = ~aif.pclk;
 
  
  
  initial begin
    uvm_config_db#(virtual apb_if)::set(null, "*", "aif", aif);
    run_test("test");
   end
endmodule
  