class sco extends uvm_scoreboard;
`uvm_component_utils(sco)

uvm_analysis_imp#(transaction , sco) recv;

bit [31:0] arr[32]= '{default:0};
bit [31:0]addr =0;
bit [31:0] data_rd=0;

function new(input string name = "sco", uvm_component parent = null);
    super.new(name,parent);
    endfunction
    
    virtual function void build_phase(uvm_phase phase);
    super.build_phase(phase);
    recv = new("recv", this);
    endfunction

virtual function void write(transaction tr);
if(tr.op == 2'd0) 
    begin 
        `uvm_info("SCO", "SYSTEM RESET DETECTED", UVM_NONE);
    end

 else if (tr.op ==2'd1)
    begin
            if(tr.pslverr == 1'b1)
                begin
                  `uvm_info("SCO", "SLV ERROR during WRITE OP", UVM_NONE);
                 end
            else 
                begin
                    arr[tr.paddr]= tr.pwdata;
                   `uvm_info("SCO", $sformatf("DATA WRITE OP  addr:%0d, wdata:%0d arr_wr:%0d",tr.paddr,tr.pwdata,  arr[tr.paddr]), UVM_NONE);
                end
     end
else if(tr.op==2'd2)
begin
            if(tr.pslverr == 1'b1)
                begin
                  `uvm_info("SCO", "SLV ERROR during WRITE OP", UVM_NONE);
                 end
            else 
                begin
                    data_rd=arr[tr.paddr];
                   //`uvm_info("SCO", $sformatf("DATA WRITE OP  addr:%0d, wdata:%0d arr_wr:%0d",tr.paddr,tr.pwdata,  arr[tr.paddr]), UVM_NONE);
                    if(data_rd == tr.prdata) begin
                      `uvm_info("SCO", $sformatf("DATA MATCHED : addr:%0d, rdata:%0d",tr.paddr,tr.prdata), UVM_NONE);end
                    else begin
                     
                      `uvm_info("SCO",$sformatf("TEST FAILED : addr:%0d, rdata:%0d data_rd_arr:%0d",tr.paddr,tr.prdata,data_rd), UVM_NONE);end
                 end

end
$display("----------------------------------------------------------------");

endfunction
 
endclass